--MATTHEW CHU
--binary2ssd.vhd
--11/7/2018
--hex display code
LIBRARY ieee;
USE ieee.STD_LOGIC_1164.all;
USE ieee.numeric_std.all;

ENTITY binary2ssd IS
	PORT (In_num    			: IN   STD_LOGIC_VECTOR(9 downto 0);
         HEX3,HEX2,HEX1,HEX0     : OUT  STD_LOGIC_VECTOR(6 downto 0));
END binary2ssd;

ARCHITECTURE behavioral of binary2ssd IS
SIGNAL thousands_dig,hundreds_dig,tens_dig,ones_dig : STD_LOGIC_VECTOR(9 DOWNTO 0);
	CONSTANT ZERO	 :STD_LOGIC_VECTOR(6 DOWNTO 0):="1000000";
	CONSTANT ONE	 :STD_LOGIC_VECTOR(6 DOWNTO 0):="1111001";
	CONSTANT TWO 	 :STD_LOGIC_VECTOR(6 DOWNTO 0):="0100100";
	CONSTANT THREE   :STD_LOGIC_VECTOR(6 DOWNTO 0):="0110000";
	CONSTANT FOUR 	 :STD_LOGIC_VECTOR(6 DOWNTO 0):="0011001";
	CONSTANT FIVE 	 :STD_LOGIC_VECTOR(6 DOWNTO 0):="0010010";
	CONSTANT SIX 	 :STD_LOGIC_VECTOR(6 DOWNTO 0):="0000010";
	CONSTANT SEVEN   :STD_LOGIC_VECTOR(6 DOWNTO 0):="1111000";
	CONSTANT EIGHT   :STD_LOGIC_VECTOR(6 DOWNTO 0):="0000000";
	CONSTANT NINE    :STD_LOGIC_VECTOR(6 DOWNTO 0):="0010000";
	CONSTANT DASH    :STD_LOGIC_VECTOR(6 DOWNTO 0):="0111111";
	CONSTANT BLANK   :STD_LOGIC_VECTOR(6 DOWNTO 0):="1111111";
BEGIN 
	--THOUSANDS
	HEX3 <= ZERO;
	--HUNDREDS
	PROCESS(In_num,hundreds_dig)
		BEGIN
			hundreds_dig <= STD_LOGIC_VECTOR(UNSIGNED(In_num)/("0001100100"));
			CASE hundreds_dig IS
				WHEN "0000000000" => HEX2 <= ZERO;
				WHEN "0000000001" => HEX2 <= ONE;
				WHEN "0000000010" => HEX2 <= TWO;
				WHEN "0000000011" => HEX2 <= THREE;
				WHEN "0000000100" => HEX2 <= FOUR;
				WHEN "0000000101" => HEX2 <= FIVE;
				WHEN "0000000110" => HEX2 <= SIX;
				WHEN "0000000111" => HEX2 <= SEVEN;
				WHEN "0000001000" => HEX2 <= EIGHT;
				WHEN "0000001001" => HEX2 <= NINE;
				WHEN OTHERS 	 => HEX2 <= BLANK;
			END CASE;
	END PROCESS;
	--TENS
	PROCESS(In_num,tens_dig)
		BEGIN
			tens_dig <= STD_LOGIC_VECTOR(UNSIGNED(In_num) rem ("0001100100")/("0000001010"));
			CASE tens_dig IS
				WHEN "0000000000" => HEX1 <= ZERO;
				WHEN "0000000001" => HEX1 <= ONE;
				WHEN "0000000010" => HEX1 <= TWO;
				WHEN "0000000011" => HEX1 <= THREE;
				WHEN "0000000100" => HEX1 <= FOUR;
				WHEN "0000000101" => HEX1 <= FIVE;
				WHEN "0000000110" => HEX1 <= SIX;
				WHEN "0000000111" => HEX1 <= SEVEN;
				WHEN "0000001000" => HEX1 <= EIGHT;
				WHEN "0000001001" => HEX1 <= NINE;
				WHEN OTHERS 	 => HEX1 <= BLANK;
			END CASE;
	END PROCESS;
	--ONES
	PROCESS(In_num,ones_dig)
		BEGIN
			ones_dig <= STD_LOGIC_VECTOR(UNSIGNED(In_num) rem ("0000001010"));
			CASE ones_dig IS
				WHEN "0000000000" => HEX0 <= ZERO;
				WHEN "0000000001" => HEX0 <= ONE;
				WHEN "0000000010" => HEX0 <= TWO;
				WHEN "0000000011" => HEX0 <= THREE;
				WHEN "0000000100" => HEX0 <= FOUR;
				WHEN "0000000101" => HEX0 <= FIVE;
				WHEN "0000000110" => HEX0 <= SIX;
				WHEN "0000000111" => HEX0 <= SEVEN;
				WHEN "0000001000" => HEX0 <= EIGHT;
				WHEN "0000001001" => HEX0 <= NINE;
				WHEN OTHERS 	 => HEX0 <= BLANK;
			END CASE;
	END PROCESS;
END behavioral;